** circuit file for profile: dff 

** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT PROFILES

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of pspice91.ini file:
.lib "D:\my_lib\orcad.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 30us 0 
.PROBE 
.INC "driver-SCHEMATIC1.net" 

.INC "driver-SCHEMATIC1.als"


.END
